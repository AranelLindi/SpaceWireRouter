----------------------------------------------------------------------------------
-- Company: University of Wuerzburg, Germany
-- Engineer: Stefan Lindoerfer
-- 
-- Create Date: 03.08.2021 20:15
-- Design Name: SpaceWire Router - Table Arbiter
-- Module Name: spwrouterarb_table
-- Project Name: Bachelor Thesis: Implementation of a SpaceWire Router on an FPGA
-- Target Devices: Xilinx FPGAs
-- Tool Versions: -/-
-- Description: Grants permission to router table and registers.
--
-- Dependencies:
-- 
-- Revision:
----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY spwrouterarb_table IS
    GENERIC (
        -- Number of SpaceWire ports.
        numports : INTEGER RANGE 1 TO 32
    );
    PORT (
        -- System clock.
        clk : IN STD_LOGIC;

        -- Synchronous reset.
        rst : IN STD_LOGIC;

        -- Requests from all ports. (Bit corresponds to port)
        request : IN STD_LOGIC_VECTOR((numports - 1) DOWNTO 0);

        -- Containts which port gets access.
        granted : OUT STD_LOGIC_VECTOR((numports - 1) DOWNTO 0)
    );
END spwrouterarb_table;

ARCHITECTURE spwrouterarb_table_arch OF spwrouterarb_table IS
    CONSTANT c_initValue : STD_LOGIC_VECTOR((numports - 1) DOWNTO 0) := (0 => '1', OTHERS => '0'); -- Initial value for arbitration algorithm

    SIGNAL s_granted : STD_LOGIC_VECTOR((numports - 1) DOWNTO 0) := c_initValue; -- Important that this signal is initialized otherwise a reset is necessary until logical addressing works as expected!
BEGIN
    -- Drive output.
    granted <= s_granted;

    -- Arbitration process.
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            IF rst = '1' THEN
                -- Synchronous reset.
                s_granted <= c_initValue;
            ELSE
                -- Check each ports (except current) wheather access is required.
                -- Method: First subsequent ones and then previous ones.
                -- Since individual, independent if-conditions are generated by for-loops,
                -- that order must be reversed to keep same priority list if-elsif-conditions would have.
                -- Example: Port4: 5..6..7..0..1..2..3 --> 1..0..7..6..5

                -- To have the right priority the order was changed in unusual order.

                Arbitration_Access : FOR i IN (numports - 1) DOWNTO 0 LOOP
                    IF (s_granted(i) = '1' AND request(i) = '0') THEN
                        pre_ports : FOR j IN (i - 1) DOWNTO 0 LOOP -- [(i-1) <= j <= 0]
                            IF (request(j) = '1') THEN
                                s_granted <= STD_LOGIC_VECTOR(to_unsigned(2 ** j, s_granted'length));
                            END IF;
                        END LOOP pre_ports;

                        -- (except current port i !)

                        seq_ports : FOR k IN (numports - 1) DOWNTO (i + 1) LOOP -- [(numports-1) <= k <= (i+1)]
                            IF (request(k) = '1') THEN
                                s_granted <= STD_LOGIC_VECTOR(to_unsigned(2 ** k, s_granted'length));
                            END IF;
                        END LOOP seq_ports;
                    END IF;
                END LOOP Arbitration_Access;
            END IF;
        END IF;
    END PROCESS;
END spwrouterarb_table_arch;